/*
inputs: sphere[4], p0[3], p1[3], BOUNDED, THRESHOLD
outputs: px0[3], px1[3], READY
*/
module ray_sphere_intersection() begin

endmodule