module scene_manager(input CLK, input MEM_READY, output[18:0] ADDRESS, output[3:0] PIXEL, output RT_READY);

/*
	this module determines what the raytracers write to in memory. 
*/

endmodule