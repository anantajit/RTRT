/*
This is a massive state machine that runs through the raytracing code. It accepts the scene data as inputs, but the mechanism for this still needs to be determined. 
*/

 module RTcore(input CLK, input[9:0] X, input[8:0] Y, output OUTPUT_READY, output[3:0] OUTPUT_PIXEL);
 
 
 
 endmodule